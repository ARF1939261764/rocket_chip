module top(

);

ChipTop ChipTop_inst();

endmodule
